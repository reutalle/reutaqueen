my_pll_inst : my_pll PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
